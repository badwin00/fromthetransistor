module hello;

initial begin
  $display("Hello World by Sam");
  $finish;
end

endmodule
